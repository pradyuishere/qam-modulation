module demodulator (
  
  );
